module pcie_x1_bfm_tb (perstn, refclkp, refclkn, hdinp0, hdinn0, hdoutp0, hdoutn0);

input wire perstn, refclkp, refclkn, hdinp0, hdinn0;
output wire hdoutp0, hdoutn0;





endmodule
